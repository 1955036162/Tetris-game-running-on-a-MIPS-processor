module test2(
    input in,
);

endmodule // 