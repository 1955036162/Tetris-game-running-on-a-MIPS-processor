module (
    
);

endmodule // 